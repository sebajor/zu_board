//default_nettype none


// This wrapper is only to simulate, the one used when compiling is generated  by vivado
module system_wrapper (
	output wire mpsoc_clk_100,
	//HPM0_FPD signals
	output wire  [39:0] HPM0_FPD_M00_axil_araddr,
	output wire  [2:0] HPM0_FPD_M00_axil_arprot,
	input wire HPM0_FPD_M00_axil_arready,
	output wire HPM0_FPD_M00_axil_arvalid,
	output wire  [39:0] HPM0_FPD_M00_axil_awaddr,
	output wire  [2:0] HPM0_FPD_M00_axil_awprot,
	input wire HPM0_FPD_M00_axil_awready,
	output wire HPM0_FPD_M00_axil_awvalid,
	output wire HPM0_FPD_M00_axil_bready,
	input wire  [1:0] HPM0_FPD_M00_axil_bresp,
	input wire HPM0_FPD_M00_axil_bvalid,
	input wire  [31:0] HPM0_FPD_M00_axil_rdata,
	output wire HPM0_FPD_M00_axil_rready,
	input wire  [1:0] HPM0_FPD_M00_axil_rresp,
	input wire HPM0_FPD_M00_axil_rvalid,
	output wire  [31:0] HPM0_FPD_M00_axil_wdata,
	input wire HPM0_FPD_M00_axil_wready,
	output wire  [3:0] HPM0_FPD_M00_axil_wstrb,
	output wire HPM0_FPD_M00_axil_wvalid,
	output wire  [39:0] HPM0_FPD_M01_axil_araddr,
	output wire  [2:0] HPM0_FPD_M01_axil_arprot,
	input wire HPM0_FPD_M01_axil_arready,
	output wire HPM0_FPD_M01_axil_arvalid,
	output wire  [39:0] HPM0_FPD_M01_axil_awaddr,
	output wire  [2:0] HPM0_FPD_M01_axil_awprot,
	input wire HPM0_FPD_M01_axil_awready,
	output wire HPM0_FPD_M01_axil_awvalid,
	output wire HPM0_FPD_M01_axil_bready,
	input wire  [1:0] HPM0_FPD_M01_axil_bresp,
	input wire HPM0_FPD_M01_axil_bvalid,
	input wire  [31:0] HPM0_FPD_M01_axil_rdata,
	output wire HPM0_FPD_M01_axil_rready,
	input wire  [1:0] HPM0_FPD_M01_axil_rresp,
	input wire HPM0_FPD_M01_axil_rvalid,
	output wire  [31:0] HPM0_FPD_M01_axil_wdata,
	input wire HPM0_FPD_M01_axil_wready,
	output wire  [3:0] HPM0_FPD_M01_axil_wstrb,
	output wire HPM0_FPD_M01_axil_wvalid,
	output wire  [39:0] HPM0_FPD_M02_axil_araddr,
	output wire  [2:0] HPM0_FPD_M02_axil_arprot,
	input wire HPM0_FPD_M02_axil_arready,
	output wire HPM0_FPD_M02_axil_arvalid,
	output wire  [39:0] HPM0_FPD_M02_axil_awaddr,
	output wire  [2:0] HPM0_FPD_M02_axil_awprot,
	input wire HPM0_FPD_M02_axil_awready,
	output wire HPM0_FPD_M02_axil_awvalid,
	output wire HPM0_FPD_M02_axil_bready,
	input wire  [1:0] HPM0_FPD_M02_axil_bresp,
	input wire HPM0_FPD_M02_axil_bvalid,
	input wire  [31:0] HPM0_FPD_M02_axil_rdata,
	output wire HPM0_FPD_M02_axil_rready,
	input wire  [1:0] HPM0_FPD_M02_axil_rresp,
	input wire HPM0_FPD_M02_axil_rvalid,
	output wire  [31:0] HPM0_FPD_M02_axil_wdata,
	input wire HPM0_FPD_M02_axil_wready,
	output wire  [3:0] HPM0_FPD_M02_axil_wstrb,
	output wire HPM0_FPD_M02_axil_wvalid,
	output wire  [39:0] HPM0_FPD_M03_axil_araddr,
	output wire  [2:0] HPM0_FPD_M03_axil_arprot,
	input wire HPM0_FPD_M03_axil_arready,
	output wire HPM0_FPD_M03_axil_arvalid,
	output wire  [39:0] HPM0_FPD_M03_axil_awaddr,
	output wire  [2:0] HPM0_FPD_M03_axil_awprot,
	input wire HPM0_FPD_M03_axil_awready,
	output wire HPM0_FPD_M03_axil_awvalid,
	output wire HPM0_FPD_M03_axil_bready,
	input wire  [1:0] HPM0_FPD_M03_axil_bresp,
	input wire HPM0_FPD_M03_axil_bvalid,
	input wire  [31:0] HPM0_FPD_M03_axil_rdata,
	output wire HPM0_FPD_M03_axil_rready,
	input wire  [1:0] HPM0_FPD_M03_axil_rresp,
	input wire HPM0_FPD_M03_axil_rvalid,
	output wire  [31:0] HPM0_FPD_M03_axil_wdata,
	input wire HPM0_FPD_M03_axil_wready,
	output wire  [3:0] HPM0_FPD_M03_axil_wstrb,
	output wire HPM0_FPD_M03_axil_wvalid,
	output wire  [39:0] HPM0_FPD_M04_axil_araddr,
	output wire  [2:0] HPM0_FPD_M04_axil_arprot,
	input wire HPM0_FPD_M04_axil_arready,
	output wire HPM0_FPD_M04_axil_arvalid,
	output wire  [39:0] HPM0_FPD_M04_axil_awaddr,
	output wire  [2:0] HPM0_FPD_M04_axil_awprot,
	input wire HPM0_FPD_M04_axil_awready,
	output wire HPM0_FPD_M04_axil_awvalid,
	output wire HPM0_FPD_M04_axil_bready,
	input wire  [1:0] HPM0_FPD_M04_axil_bresp,
	input wire HPM0_FPD_M04_axil_bvalid,
	input wire  [31:0] HPM0_FPD_M04_axil_rdata,
	output wire HPM0_FPD_M04_axil_rready,
	input wire  [1:0] HPM0_FPD_M04_axil_rresp,
	input wire HPM0_FPD_M04_axil_rvalid,
	output wire  [31:0] HPM0_FPD_M04_axil_wdata,
	input wire HPM0_FPD_M04_axil_wready,
	output wire  [3:0] HPM0_FPD_M04_axil_wstrb,
	output wire HPM0_FPD_M04_axil_wvalid,
	output wire axil_arst_n, axil_rst
);



endmodule
`resetall